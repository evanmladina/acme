library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.Types.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(-432);
    constant feature : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 0, 0, 0, -2, -2, 3, -2, -2, 3, 4, -2, -2, 0, -2, -2, 3, 4, 0, -2, -2, 3, -2, -2, 3, 2, -2, -2, 4, -2, -2),
                (0, 0, 0, 0, -2, -2, 3, -2, -2, 3, 4, -2, -2, 0, -2, -2, 0, 3, 4, -2, -2, 4, -2, -2, 4, 0, -2, -2, 3, -2, -2),
                (0, 0, 0, 0, -2, -2, 3, -2, -2, 3, 2, -2, -2, 0, -2, -2, 0, 3, 4, -2, -2, 4, -2, -2, 4, 0, -2, -2, 3, -2, -2),
                (0, 0, 0, -2, 0, -2, -2, 0, 3, -2, -2, 4, -2, -2, 0, 4, 1, -2, -2, 3, -2, -2, 4, 0, -2, -2, 3, -2, -2, -2, -2),
                (0, 0, 0, 0, -2, -2, 3, -2, -2, 3, 0, -2, -2, 1, -2, -2, 0, 4, 0, -2, -2, 3, -2, -2, 4, 0, -2, -2, 3, -2, -2),
                (0, 0, 0, -2, 0, -2, -2, 3, 2, -2, -2, 1, -2, -2, 0, 4, 1, -2, -2, 3, -2, -2, 4, 0, -2, -2, 3, -2, -2, -2, -2),
                (0, 0, 0, -2, 0, -2, -2, 3, 1, -2, -2, 1, -2, -2, 0, 4, 3, -2, -2, 3, -2, -2, 4, 0, -2, -2, 3, -2, -2, -2, -2),
                (0, 0, 0, -2, 3, -2, -2, 3, 4, -2, -2, 1, -2, -2, 0, 4, 3, -2, -2, 3, -2, -2, 4, 0, -2, -2, 3, -2, -2, -2, -2),
                (0, 0, 0, -2, 0, -2, -2, 3, 2, -2, -2, 0, -2, -2, 0, 3, 2, -2, -2, 2, -2, -2, 4, 0, -2, -2, 0, -2, -2, -2, -2),
                (0, 0, 0, -2, 4, -2, -2, 1, 1, -2, -2, 0, -2, -2, 0, 4, 0, -2, -2, 3, -2, -2, 4, 0, -2, -2, 0, -2, -2, -2, -2),
                (0, 0, 0, 0, -2, -2, 4, -2, -2, 1, 4, -2, -2, 3, -2, -2, 0, 4, 1, -2, -2, 3, -2, -2, 4, 0, -2, -2, 3, -2, -2),
                (0, 0, 4, 0, -2, -2, 3, -2, -2, 3, 2, -2, -2, 2, -2, -2, 0, 1, 1, -2, -2, 3, -2, -2, 4, 0, -2, -2, 0, -2, -2),
                (0, 0, 0, 4, -2, -2, 4, -2, -2, 1, 1, -2, -2, 4, -2, -2, 0, 4, 1, -2, -2, 2, -2, -2, 4, 0, -2, -2, 3, -2, -2),
                (0, 3, 0, 0, -2, -2, 4, -2, -2, 1, 3, -2, -2, 2, -2, -2, 0, 4, 1, -2, -2, 3, -2, -2, 4, 1, -2, -2, 2, -2, -2),
                (0, 3, 2, 1, -2, -2, 3, -2, -2, 3, 2, -2, -2, 1, -2, -2, 0, 4, 0, -2, -2, 3, -2, -2, 4, 0, -2, -2, 0, -2, -2),
                (0, 0, 3, 1, -2, -2, 0, -2, -2, 1, 1, -2, -2, 3, -2, -2, 0, 1, 1, -2, -2, 3, -2, -2, 2, 4, -2, -2, 3, -2, -2),
                (0, 0, 0, 4, -2, -2, 4, -2, -2, 2, 4, -2, -2, 1, -2, -2, 0, 4, 1, -2, -2, 2, -2, -2, 4, 3, -2, -2, 0, -2, -2),
                (0, 0, 3, 2, -2, -2, 1, -2, -2, 4, 1, -2, -2, 2, -2, -2, 4, 3, 0, -2, -2, 0, -2, -2, 3, 2, -2, -2, 2, -2, -2),
                (0, 0, 0, 0, -2, -2, 4, -2, -2, 4, 1, -2, -2, 2, -2, -2, 3, 2, 3, -2, -2, 3, -2, -2, 4, 3, -2, -2, 0, -2, -2),
                (0, 0, 3, 2, -2, -2, 1, -2, -2, 1, 1, -2, -2, 3, -2, -2, 4, 3, 0, -2, -2, 0, -2, -2, 3, 2, -2, -2, 2, -2, -2),
                (0, 0, 0, 0, -2, -2, 4, -2, -2, 2, 3, -2, -2, 2, -2, -2, 3, 0, 3, -2, -2, 2, -2, -2, 4, 0, -2, -2, 2, -2, -2),
                (0, 0, 3, 1, -2, -2, 1, -2, -2, 2, 3, -2, -2, 3, -2, -2, 4, 3, 0, -2, -2, 2, -2, -2, 3, 2, -2, -2, 2, -2, -2),
                (0, 0, 3, 2, -2, -2, 1, -2, -2, 1, 1, -2, -2, 0, -2, -2, 3, 0, 2, -2, -2, 2, -2, -2, 0, 0, -2, -2, 3, -2, -2),
                (3, 0, 0, 3, -2, -2, 1, -2, -2, 2, 3, -2, -2, 0, -2, -2, 0, 2, 1, -2, -2, 1, -2, -2, 0, 2, -2, -2, 3, -2, -2),
                (3, 0, 3, 2, -2, -2, 2, -2, -2, 2, 3, -2, -2, 0, -2, -2, 3, 0, 2, -2, -2, 4, -2, -2, 4, 3, -2, -2, 0, -2, -2),
                (3, 0, 0, 2, -2, -2, 1, -2, -2, 2, 3, -2, -2, 0, -2, -2, 3, 2, 0, -2, -2, 0, -2, -2, 0, 3, -2, -2, 3, -2, -2),
                (3, 0, 0, 0, -2, -2, 1, -2, -2, 2, 1, -2, -2, 0, -2, -2, 3, 0, 2, -2, -2, 4, -2, -2, 0, 3, -2, -2, 3, -2, -2),
                (3, 2, 0, 1, -2, -2, 1, -2, -2, 3, 0, -2, -2, 2, -2, -2, 3, 2, 0, -2, -2, 0, -2, -2, 0, 0, -2, -2, 3, -2, -2),
                (3, 2, 0, 1, -2, -2, 3, -2, -2, 3, 0, -2, -2, 2, -2, -2, 2, 0, 4, -2, -2, 4, -2, -2, 3, 0, -2, -2, 1, -2, -2),
                (3, 2, 4, 0, -2, -2, 3, -2, -2, 0, 0, -2, -2, 3, -2, -2, 2, 0, 1, -2, -2, 2, -2, -2, 3, 0, -2, -2, 0, -2, -2),
                (3, 0, 4, 1, -2, -2, 3, -2, -2, 2, 3, -2, -2, 0, -2, -2, 2, 2, 0, -2, -2, 3, -2, -2, 4, 1, -2, -2, 0, -2, -2),
                (3, 2, 3, 0, -2, -2, 4, -2, -2, 0, 3, -2, -2, 1, -2, -2, 2, 1, 2, -2, -2, 1, -2, -2, 3, 0, -2, -2, 1, -2, -2),
                (3, 1, 0, 4, -2, -2, 2, -2, -2, 1, 0, -2, -2, 0, -2, -2, 2, 0, 1, -2, -2, 4, -2, -2, 2, 3, -2, -2, 0, -2, -2),
                (3, 0, 0, 3, -2, -2, 4, -2, -2, 1, 1, -2, -2, 0, -2, -2, 0, 0, 3, -2, -2, 4, -2, -2, 3, 4, -2, -2, 4, -2, -2),
                (3, 2, 3, 0, -2, -2, 4, -2, -2, 0, 4, -2, -2, 0, -2, -2, 2, 0, 2, -2, -2, 3, -2, -2, 1, 4, -2, -2, 4, -2, -2),
                (3, 0, 0, 0, -2, -2, 2, -2, -2, 2, 0, -2, -2, 4, -2, -2, 2, 1, 2, -2, -2, 1, -2, -2, 2, 3, -2, -2, 0, -2, -2),
                (3, 2, 4, 1, -2, -2, 2, -2, -2, 0, 1, -2, -2, 4, -2, -2, 2, 1, 2, -2, -2, 1, -2, -2, 1, 1, -2, -2, 1, -2, -2),
                (3, 0, 0, 2, -2, -2, 1, -2, -2, 2, 4, -2, -2, 3, -2, -2, 2, 4, 0, -2, -2, 2, -2, -2, 2, 1, -2, -2, 2, -2, -2),
                (0, 0, 3, 2, -2, -2, 4, -2, -2, 0, 3, -2, -2, 4, -2, -2, 1, 1, 4, -2, -2, 2, -2, -2, 0, 0, -2, -2, 2, -2, -2),
                (3, 2, 0, 1, -2, -2, 0, -2, -2, 0, 2, -2, -2, 2, -2, -2, 2, 4, 0, -2, -2, 2, -2, -2, 2, 1, -2, -2, 3, -2, -2),
                (3, 0, 0, 2, -2, -2, 2, -2, -2, 2, 4, -2, -2, 2, -2, -2, 2, 4, 1, -2, -2, 2, -2, -2, 2, 1, -2, -2, 2, -2, -2),
                (3, 0, 4, 1, -2, -2, 2, -2, -2, 4, 2, -2, -2, 3, -2, -2, 0, 0, 4, -2, -2, 3, -2, -2, 4, 0, -2, -2, 3, -2, -2),
                (0, 0, 3, 2, -2, -2, 4, -2, -2, 2, 1, -2, -2, 2, -2, -2, 1, 1, 3, -2, -2, 2, -2, -2, 4, 0, -2, -2, 4, -2, -2),
                (3, 2, 0, 1, -2, -2, 3, -2, -2, 0, 2, -2, -2, 2, -2, -2, 2, 4, 0, -2, -2, 1, -2, -2, 2, 4, -2, -2, 0, -2, -2),
                (3, 0, 4, 0, -2, -2, 2, -2, -2, 4, 3, -2, -2, 3, -2, -2, 0, 2, 0, -2, -2, 0, -2, -2, 0, 1, -2, -2, 4, -2, -2),
                (1, 3, 0, 4, -2, -2, 2, -2, -2, 2, 0, -2, -2, 2, -2, -2, 1, 0, 0, -2, -2, 2, -2, -2, 4, 0, -2, -2, 0, -2, -2),
                (0, 0, 3, 2, -2, -2, 4, -2, -2, 1, 3, -2, -2, 1, -2, -2, 1, 1, 4, -2, -2, 2, -2, -2, 3, 2, -2, -2, 4, -2, -2),
                (2, 0, 4, 0, -2, -2, 0, -2, -2, 4, 3, -2, -2, 3, -2, -2, 0, 4, 1, -2, -2, 0, -2, -2, 2, 3, -2, -2, 2, -2, -2),
                (3, 0, 0, 0, -2, -2, 3, -2, -2, 2, 3, -2, -2, 3, -2, -2, 0, 0, 0, -2, -2, 4, -2, -2, 3, 4, -2, -2, 4, -2, -2),
                (3, 0, 0, 2, -2, -2, 2, -2, -2, 2, 4, -2, -2, 4, -2, -2, 2, 4, 1, -2, -2, 1, -2, -2, 2, 4, -2, -2, 2, -2, -2),
                (1, 3, 0, 4, -2, -2, 2, -2, -2, 2, 0, -2, -2, 2, -2, -2, 1, 0, 0, -2, -2, 2, -2, -2, 3, 0, -2, -2, 3, -2, -2),
                (0, 0, 0, 0, -2, -2, 1, -2, -2, 3, 2, -2, -2, 3, -2, -2, 0, 3, 3, -2, -2, 4, -2, -2, 4, 1, -2, -2, 3, -2, -2),
                (3, 0, 4, 0, -2, -2, 0, -2, -2, 4, 3, -2, -2, 4, -2, -2, 0, 0, 3, -2, -2, 3, -2, -2, 3, 4, -2, -2, 4, -2, -2),
                (1, 4, 3, 0, -2, -2, 0, -2, -2, 0, 3, -2, -2, 3, -2, -2, 1, 1, 0, -2, -2, 0, -2, -2, 4, 0, -2, -2, 4, -2, -2),
                (3, 0, 4, 0, -2, -2, 2, -2, -2, 4, 0, -2, -2, 3, -2, -2, 4, 0, 3, -2, -2, 4, -2, -2, 0, 4, -2, -2, 4, -2, -2),
                (3, 0, 0, 2, -2, -2, 2, -2, -2, 2, 4, -2, -2, 0, -2, -2, 2, 4, 0, -2, -2, 2, -2, -2, 0, 0, -2, -2, 3, -2, -2),
                (2, 2, 4, 3, -2, -2, 0, -2, -2, 0, 3, -2, -2, 1, -2, -2, 0, 0, 0, -2, -2, 0, -2, -2, 3, 0, -2, -2, 4, -2, -2),
                (1, 1, 3, 0, -2, -2, 4, -2, -2, 1, 1, -2, -2, 3, -2, -2, 0, 0, 4, -2, -2, 4, -2, -2, 4, 4, -2, -2, 4, -2, -2),
                (0, 0, 0, 0, -2, -2, 2, -2, -2, 3, 2, -2, -2, 1, -2, -2, 0, 3, 4, -2, -2, 4, -2, -2, 4, 1, -2, -2, 3, -2, -2),
                (2, 4, 3, 0, -2, -2, 2, -2, -2, 0, 2, -2, -2, 2, -2, -2, 0, 4, 0, -2, -2, 3, -2, -2, 3, 2, -2, -2, 0, -2, -2),
                (3, 0, 4, 0, -2, -2, 2, -2, -2, 2, 0, -2, -2, 2, -2, -2, 0, 0, 2, -2, -2, 4, -2, -2, 4, 0, -2, -2, 2, -2, -2),
                (1, 4, 3, 0, -2, -2, 4, -2, -2, 0, 2, -2, -2, 3, -2, -2, 1, 1, 4, -2, -2, 4, -2, -2, 4, 0, -2, -2, 4, -2, -2),
                (2, 3, 0, 4, -2, -2, 2, -2, -2, 0, 4, -2, -2, 4, -2, -2, 0, 2, 3, -2, -2, 0, -2, -2, 1, 1, -2, -2, 4, -2, -2),
                (1, 1, 3, 0, -2, -2, 3, -2, -2, 1, 1, -2, -2, 2, -2, -2, 0, 0, 4, -2, -2, 4, -2, -2, 4, 4, -2, -2, 4, -2, -2),
                (3, 0, 0, 0, -2, -2, 2, -2, -2, 2, 4, -2, -2, 1, -2, -2, 2, 4, 0, -2, -2, 2, -2, -2, 2, 4, -2, -2, 0, -2, -2),
                (0, 0, 4, 2, -2, -2, 2, -2, -2, 3, 2, -2, -2, 3, -2, -2, 3, 2, 4, -2, -2, 4, -2, -2, 2, 0, -2, -2, 1, -2, -2),
                (3, 0, 4, 0, -2, -2, 2, -2, -2, 2, 0, -2, -2, 3, -2, -2, 0, 3, 1, -2, -2, 0, -2, -2, 4, 3, -2, -2, 1, -2, -2),
                (3, 0, 4, 0, -2, -2, 0, -2, -2, 4, 3, -2, -2, 2, -2, -2, 4, 0, 0, -2, -2, 3, -2, -2, 2, 4, -2, -2, 3, -2, -2),
                (3, 0, 2, 3, -2, -2, 0, -2, -2, 2, 4, -2, -2, 4, -2, -2, 2, 4, 0, -2, -2, 2, -2, -2, 2, 0, -2, -2, 0, -2, -2),
                (3, 0, 4, 1, -2, -2, 1, -2, -2, 2, 3, -2, -2, 3, -2, -2, 2, 0, 0, -2, -2, 4, -2, -2, 1, 0, -2, -2, 1, -2, -2),
                (3, 0, 4, 0, -2, -2, 2, -2, -2, 2, 0, -2, -2, 2, -2, -2, 0, 0, 1, -2, -2, 1, -2, -2, 4, 3, -2, -2, 3, -2, -2),
                (3, 0, 4, 0, -2, -2, 2, -2, -2, 2, 4, -2, -2, 3, -2, -2, 0, 3, 1, -2, -2, 0, -2, -2, 4, 3, -2, -2, 1, -2, -2),
                (2, 2, 4, 3, -2, -2, 1, -2, -2, 0, 3, -2, -2, 1, -2, -2, 0, 4, 1, -2, -2, 0, -2, -2, 3, 2, -2, -2, 4, -2, -2),
                (1, 0, 0, 2, -2, -2, 1, -2, -2, 2, 2, -2, -2, 1, -2, -2, 0, 4, 3, -2, -2, 4, -2, -2, 4, 4, -2, -2, 0, -2, -2),
                (3, 0, 4, 2, -2, -2, 2, -2, -2, 2, 3, -2, -2, 3, -2, -2, 0, 3, 1, -2, -2, 0, -2, -2, 0, 4, -2, -2, 3, -2, -2),
                (0, 4, 3, 0, -2, -2, 0, -2, -2, 1, 0, -2, -2, 2, -2, -2, 3, 4, 0, -2, -2, 3, -2, -2, 3, 4, -2, -2, 2, -2, -2),
                (1, 1, 3, 0, -2, -2, 2, -2, -2, 1, 1, -2, -2, 3, -2, -2, 0, 0, 4, -2, -2, 2, -2, -2, 4, 4, -2, -2, 2, -2, -2),
                (2, 4, 3, 0, -2, -2, 2, -2, -2, 0, 2, -2, -2, 2, -2, -2, 0, 4, 0, -2, -2, 2, -2, -2, 3, 3, -2, -2, 4, -2, -2),
                (0, 0, 4, 1, -2, -2, 2, -2, -2, 1, 1, -2, -2, 4, -2, -2, 3, 2, 4, -2, -2, 0, -2, -2, 1, 2, -2, -2, 4, -2, -2),
                (3, 0, 2, 3, -2, -2, 0, -2, -2, 2, 4, -2, -2, 4, -2, -2, 2, 4, 2, -2, -2, 0, -2, -2, 0, 1, -2, -2, 1, -2, -2),
                (3, 0, 4, 1, -2, -2, 3, -2, -2, 2, 0, -2, -2, 4, -2, -2, 2, 0, 0, -2, -2, 4, -2, -2, 1, 4, -2, -2, 1, -2, -2),
                (1, 2, 4, 0, -2, -2, 2, -2, -2, 0, 4, -2, -2, 3, -2, -2, 4, 0, 4, -2, -2, 4, -2, -2, 0, 2, -2, -2, 2, -2, -2),
                (3, 0, 4, 3, -2, -2, 2, -2, -2, 2, 2, -2, -2, 0, -2, -2, 2, 1, 3, -2, -2, 0, -2, -2, 1, 0, -2, -2, 1, -2, -2),
                (3, 0, 4, 0, -2, -2, 2, -2, -2, 2, 2, -2, -2, 3, -2, -2, 2, 0, 0, -2, -2, 0, -2, -2, 1, 0, -2, -2, 0, -2, -2),
                (0, 4, 2, 4, -2, -2, 0, -2, -2, 2, 0, -2, -2, 3, -2, -2, 3, 4, 4, -2, -2, 0, -2, -2, 2, 2, -2, -2, 3, -2, -2),
                (3, 0, 4, 0, -2, -2, 2, -2, -2, 4, 2, -2, -2, 2, -2, -2, 1, 0, 1, -2, -2, 0, -2, -2, 3, 4, -2, -2, 3, -2, -2),
                (2, 2, 3, 0, -2, -2, 2, -2, -2, 0, 4, -2, -2, 1, -2, -2, 1, 1, 2, -2, -2, 3, -2, -2, 4, 1, -2, -2, 1, -2, -2),
                (3, 0, 4, 0, -2, -2, 1, -2, -2, 2, 2, -2, -2, 4, -2, -2, 3, 2, 4, -2, -2, 1, -2, -2, 3, 2, -2, -2, 2, -2, -2),
                (1, 2, 4, 0, -2, -2, 2, -2, -2, 0, 4, -2, -2, 3, -2, -2, 0, 4, 3, -2, -2, 4, -2, -2, 4, 4, -2, -2, 2, -2, -2),
                (3, 0, 2, 3, -2, -2, 0, -2, -2, 2, 4, -2, -2, 0, -2, -2, 2, 4, 0, -2, -2, 4, -2, -2, 0, 1, -2, -2, 1, -2, -2),
                (3, 0, 4, 1, -2, -2, 1, -2, -2, 2, 3, -2, -2, 4, -2, -2, 2, 0, 1, -2, -2, 2, -2, -2, 1, 0, -2, -2, 1, -2, -2),
                (3, 0, 4, 4, -2, -2, 2, -2, -2, 4, 4, -2, -2, 2, -2, -2, 0, 2, 0, -2, -2, 2, -2, -2, 2, 3, -2, -2, 2, -2, -2),
                (3, 0, 4, 0, -2, -2, 2, -2, -2, 2, 2, -2, -2, 0, -2, -2, 2, 4, 2, -2, -2, 3, -2, -2, 1, 2, -2, -2, 1, -2, -2),
                (1, 1, 3, 0, -2, -2, 4, -2, -2, 3, 0, -2, -2, 0, -2, -2, 4, 0, 1, -2, -2, 0, -2, -2, 4, 0, -2, -2, 2, -2, -2),
                (3, 0, 4, 4, -2, -2, 1, -2, -2, 2, 0, -2, -2, 1, -2, -2, 2, 2, 3, -2, -2, 4, -2, -2, 1, 4, -2, -2, 1, -2, -2),
                (2, 2, 4, 3, -2, -2, 1, -2, -2, 0, 4, -2, -2, 1, -2, -2, 1, 1, 3, -2, -2, 3, -2, -2, 4, 1, -2, -2, 1, -2, -2),
                (3, 0, 4, 0, -2, -2, 2, -2, -2, 2, 4, -2, -2, 4, -2, -2, 0, 4, 0, -2, -2, 2, -2, -2, 4, 3, -2, -2, 4, -2, -2),
                (0, 4, 0, 4, -2, -2, 2, -2, -2, 3, 2, -2, -2, 2, -2, -2, 3, 4, 3, -2, -2, 2, -2, -2, 2, 2, -2, -2, 0, -2, -2),
                (3, 0, 2, 4, -2, -2, 0, -2, -2, 2, 4, -2, -2, 0, -2, -2, 2, 1, 1, -2, -2, 4, -2, -2, 1, 2, -2, -2, 2, -2, -2),
                (3, 0, 1, 4, -2, -2, 1, -2, -2, 2, 4, -2, -2, 3, -2, -2, 2, 0, 4, -2, -2, 3, -2, -2, 1, 2, -2, -2, 1, -2, -2)
                );
    constant threshold_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((221, 103, 40, -66, -256, -256, 108, -256, -256, 226, -107, -256, -256, 167, -256, -256, 391, -6, 351, -256, -256, 189, -256, -256, 666, 80, -256, -256, 808, -256, -256),
                (187, 83, 26, -66, -256, -256, 61, -256, -256, 110, -107, -256, -256, 134, -256, -256, 360, 223, -87, -256, -256, -6, -256, -256, 177, 524, -256, -256, 263, -256, -256),
                (187, 76, 12, -66, -256, -256, 105, -256, -256, 83, -187, -256, -256, 137, -256, -256, 338, 223, -26, -256, -256, -6, -256, -256, 157, 465, -256, -256, 263, -256, -256),
                (181, 70, -66, -256, 2, -256, -256, 128, 66, -256, -256, -26, -256, -256, 307, -26, 127, -256, -256, 108, -256, -256, 157, 456, -256, -256, 263, -256, -256, -256, -256),
                (181, 70, 3, -66, -256, -256, 66, -256, -256, 167, 147, -256, -256, 109, -256, -256, 307, -107, 245, -256, -256, 108, -256, -256, 157, 465, -256, -256, 263, -256, -256),
                (171, 55, -66, -256, -8, -256, -256, 66, -71, -256, -256, 109, -256, -256, 307, 25, 127, -256, -256, 90, -256, -256, 177, 465, -256, -256, 263, -256, -256, -256, -256),
                (171, 65, -66, -256, 22, -256, -256, 194, 127, -256, -256, 91, -256, -256, 305, -107, 24, -256, -256, 90, -256, -256, 177, 456, -256, -256, 263, -256, -256, -256, -256),
                (164, 55, -66, -256, 56, -256, -256, 152, -107, -256, -256, 109, -256, -256, 302, -107, 12, -256, -256, 90, -256, -256, 157, 524, -256, -256, 263, -256, -256, -256, -256),
                (164, 55, -66, -256, -16, -256, -256, 68, -187, -256, -256, 111, -256, -256, 386, 108, -39, -256, -256, -9, -256, -256, 208, 544, -256, -256, 1067, -256, -256, -256, -256),
                (163, 43, -66, -256, -107, -256, -256, 109, 1, -256, -256, 144, -256, -256, 386, -107, 252, -256, -256, 81, -256, -256, 208, 571, -256, -256, 954, -256, -256, -256, -256),
                (163, 90, 5, -66, -256, -256, -107, -256, -256, 127, -57, -256, -256, 17, -256, -256, 302, 25, 109, -256, -256, 73, -256, -256, 65, 494, -256, -256, 263, -256, -256),
                (163, 38, -107, -68, -256, -256, 31, -256, -256, 31, -134, -256, -256, -35, -256, -256, 386, 109, 1, -256, -256, 17, -256, -256, 309, 524, -256, -256, 954, -256, -256),
                (147, 27, -66, -107, -256, -256, -107, -256, -256, 109, 1, -256, -256, -107, -256, -256, 302, -26, 109, -256, -256, -10, -256, -256, 177, 544, -256, -256, 263, -256, -256),
                (147, 152, -2, -66, -256, -256, -107, -256, -256, 91, 373, -256, -256, 18, -256, -256, 302, -36, 109, -256, -256, 56, -256, -256, 65, 109, -256, -256, -141, -256, -256),
                (147, 83, -228, 164, -256, -256, 12, -256, -256, 250, -7, -256, -256, 91, -256, -256, 404, -107, 245, -256, -256, 68, -256, -256, 330, 524, -256, -256, 954, -256, -256),
                (147, 26, -87, 127, -256, -256, -27, -256, -256, 109, 1, -256, -256, -28, -256, -256, 404, 109, 1, -256, -256, 4, -256, -256, -103, -6, -256, -256, 130, -256, -256),
                (145, 26, -66, -107, -256, -256, -107, -256, -256, 316, -107, -256, -256, 91, -256, -256, 390, 25, 127, -256, -256, 4, -256, -256, 309, 78, -256, -256, 1069, -256, -256),
                (275, 110, 61, -246, -256, -256, 91, -256, -256, -26, 109, -256, -256, 312, -256, -256, -107, -92, 352, -256, -256, 277, -256, -256, 93, -32, -256, -256, -44, -256, -256),
                (275, 110, -4, -66, -256, -256, -107, -256, -256, -26, 109, -256, -256, -15, -256, -256, 1072, -39, 53, -256, -256, 240, -256, -256, 2420, 2051, -256, -256, 2272, -256, -256),
                (275, 110, 31, -175, -256, -256, 109, -256, -256, 127, -35, -256, -256, -3, -256, -256, -107, -92, 352, -256, -256, 277, -256, -256, 90, -121, -256, -256, -44, -256, -256),
                (278, 90, -19, -66, -256, -256, -107, -256, -256, 25, 12, -256, -256, 312, -256, -256, 1047, 1067, 277, -256, -256, -143, -256, -256, 2420, 353, -256, -256, 291, -256, -256),
                (278, 90, 115, -53, -256, -256, 91, -256, -256, -15, 17, -256, -256, 68, -256, -256, -107, -87, 432, -256, -256, -182, -256, -256, 56, -121, -256, -256, -102, -256, -256),
                (278, 38, 110, -277, -256, -256, 109, -256, -256, 109, 37, -256, -256, 223, -256, -256, 937, 1067, 6, -256, -256, -126, -256, -256, 1971, 704, -256, -256, 2233, -256, -256),
                (250, 126, -13, -87, -256, -256, -53, -256, -256, 52, 56, -256, -256, 387, -256, -256, 340, 28, -125, -256, -256, 91, -256, -256, 956, 22, -256, -256, 833, -256, -256),
                (295, 127, 12, -162, -256, -256, -43, -256, -256, -11, 41, -256, -256, 702, -256, -256, 1072, 1282, 112, -256, -256, 309, -256, -256, 1469, 2051, -256, -256, 1235, -256, -256),
                (250, 126, 2, -277, -256, -256, 109, -256, -256, -39, 19, -256, -256, 600, -256, -256, 494, 65, 850, -256, -256, 698, -256, -256, 1492, 1072, -256, -256, 1774, -256, -256),
                (295, 127, -19, -66, -256, -256, -53, -256, -256, 55, -53, -256, -256, 627, -256, -256, 1077, 953, 117, -256, -256, 309, -256, -256, 2917, 2600, -256, -256, 2697, -256, -256),
                (250, -246, 158, 164, -256, -256, 109, -256, -256, 26, 221, -256, -256, -106, -256, -256, 494, 65, 826, -256, -256, 694, -256, -256, 1492, 464, -256, -256, 1785, -256, -256),
                (250, -282, 160, 164, -256, -256, -92, -256, -256, 56, 221, -256, -256, -39, -256, -256, 22, 822, 147, -256, -256, 157, -256, -256, 491, 751, -256, -256, -35, -256, -256),
                (149, -217, -6, 554, -256, -256, -3, -256, -256, 222, 163, -256, -256, -3, -256, -256, 24, 822, -89, -256, -256, -124, -256, -256, 494, 751, -256, -256, 221, -256, -256),
                (285, 16, -107, 1, -256, -256, -1, -256, -256, -69, 4, -256, -256, 659, -256, -256, 366, 117, 850, -256, -256, 1077, -256, -256, 86, -35, -256, -256, 121, -256, -256),
                (115, -159, -25, 553, -256, -256, -6, -256, -256, 222, -1, -256, -256, -17, -256, -256, 37, -53, -72, -256, -256, 145, -256, -256, 509, 700, -256, -256, -125, -256, -256),
                (120, -53, 219, 330, -256, -256, -171, -256, -256, 109, 63, -256, -256, 223, -256, -256, 24, 822, -89, -256, -256, 309, -256, -256, 322, 885, -256, -256, 4, -256, -256),
                (314, 2, -66, -87, -256, -256, -107, -256, -256, 127, -17, -256, -256, 223, -256, -256, 1492, 364, 676, -256, -256, 25, -256, -256, 1785, 279, -256, -256, 1337, -256, -256),
                (314, -110, 7, 596, -256, -256, -6, -256, -256, 705, 747, -256, -256, 887, -256, -256, 366, 1492, 136, -256, -256, 907, -256, -256, -17, 508, -256, -256, -46, -256, -256),
                (90, 221, 60, -29, -256, -256, -23, -256, -256, -264, 238, -256, -256, -16, -256, -256, -3, -35, -108, -256, -256, 145, -256, -256, 301, 885, -256, -256, 6, -256, -256),
                (68, -207, -6, 164, -256, -256, -222, -256, -256, 221, -53, -256, -256, -16, -256, -256, -20, -107, -150, -256, -256, 145, -256, -256, 91, 55, -256, -256, 164, -256, -256),
                (31, 653, 221, -111, -256, -256, 127, -256, -256, -217, 4, -256, -256, -11, -256, -256, -74, -6, 340, -256, -256, -159, -256, -256, 38, -53, -256, -256, 291, -256, -256),
                (2, -66, -84, -273, -256, -256, -107, -256, -256, -37, -87, -256, -256, -107, -256, -256, 109, 55, -57, -256, -256, -84, -256, -256, 544, 223, -256, -256, -172, -256, -256),
                (12, -282, 258, 164, -256, -256, 270, -256, -256, 221, -97, -256, -256, -244, -256, -256, -110, -6, 339, -256, -256, -159, -256, -256, -20, -17, -256, -256, 509, -256, -256),
                (4, 653, 221, -132, -256, -256, -245, -256, -256, -217, 4, -256, -256, -215, -256, -256, -110, -6, 145, -256, -256, -159, -256, -256, -21, -17, -256, -256, 321, -256, -256),
                (961, 937, 747, 109, -256, -256, 111, -256, -256, 137, -211, -256, -256, 622, -256, -256, 1971, 553, -107, -256, -256, 2594, -256, -256, 1337, 1977, -256, -256, 2688, -256, -256),
                (-16, -66, -84, -273, -256, -256, -107, -256, -256, -278, 73, -256, -256, 306, -256, -256, 109, 1, 314, -256, -256, -39, -256, -256, -107, 242, -256, -256, -16, -256, -256),
                (-25, -282, 258, 164, -256, -256, -87, -256, -256, 221, -181, -256, -256, -239, -256, -256, -159, -6, 338, -256, -256, 182, -256, -256, -63, 126, -256, -256, 1069, -256, -256),
                (937, 937, 777, 221, -256, -256, 111, -256, -256, 137, 917, -256, -256, 622, -256, -256, 553, 161, 512, -256, -256, 551, -256, -256, 1971, 182, -256, -256, 899, -256, -256),
                (-53, 314, 219, 330, -256, -256, -171, -256, -256, 163, 1015, -256, -256, 358, -256, -256, 109, -2, -36, -256, -256, 38, -256, -256, -107, 242, -256, -256, 223, -256, -256),
                (-23, -66, -84, -273, -256, -256, -107, -256, -256, -17, 370, -256, -256, 91, -256, -256, 109, 1, -57, -256, -256, -96, -256, -256, 1284, 146, -256, -256, 3778, -256, -256),
                (349, 1272, 747, 221, -256, -256, 849, -256, -256, 472, 1450, -256, -256, 905, -256, -256, -13, 289, 73, -256, -256, -23, -256, -256, 349, 333, -256, -256, 376, -256, -256),
                (494, 221, 205, -3, -256, -256, 420, -256, -256, 146, 108, -256, -256, 233, -256, -256, 1538, 350, 221, -256, -256, 25, -256, -256, 1785, 309, -256, -256, 1337, -256, -256),
                (-25, 506, 221, -187, -256, -256, -263, -256, -256, -200, 4, -256, -256, -6, -256, -256, -165, -16, 145, -256, -256, 218, -256, -256, -39, 147, -256, -256, 301, -256, -256),
                (-35, 250, 219, 330, -256, -256, -200, -256, -256, 250, 1649, -256, -256, 377, -256, -256, 109, -16, -47, -256, -256, 87, -256, -256, -87, 243, -256, -256, 511, -256, -256),
                (221, 205, -16, -66, -256, -256, 109, -256, -256, 420, 106, -256, -256, 427, -256, -256, 257, 705, -47, -256, -256, 15, -256, -256, -107, 164, -256, -256, 108, -256, -256),
                (1284, 1340, 747, 221, -256, -256, 849, -256, -256, 289, 265, -256, -256, 3864, -256, -256, 2917, 747, 1313, -256, -256, 2600, -256, -256, 2697, 630, -256, -256, 3259, -256, -256),
                (-35, 665, 494, 220, -256, -256, 224, -256, -256, 1071, 698, -256, -256, 771, -256, -256, 91, 73, 834, -256, -256, -2, -256, -256, -97, 242, -256, -256, -16, -256, -256),
                (1072, 891, 787, 221, -256, -256, 143, -256, -256, 65, 908, -256, -256, 622, -256, -256, 1469, 376, 1138, -256, -256, 1418, -256, -256, 1235, 1484, -256, -256, 1571, -256, -256),
                (-25, 653, 221, -128, -256, -256, -201, -256, -256, -240, 4, -256, -256, 776, -256, -256, -110, -16, 338, -256, -256, -162, -256, -256, 220, 205, -256, -256, 83, -256, -256),
                (366, 5, 147, -30, -256, -256, 682, -256, -256, 75, 152, -256, -256, 164, -256, -256, -4, -27, -66, -256, -256, -26, -256, -256, 671, 194, -256, -256, 86, -256, -256),
                (218, -35, 250, 219, -256, -256, -57, -256, -256, 91, 73, -256, -256, -84, -256, -256, 207, 207, 1204, -256, -256, 208, -256, -256, -77, -118, -256, -256, -36, -256, -256),
                (221, 205, -29, -66, -256, -256, 291, -256, -256, 420, 106, -256, -256, -53, -256, -256, 257, 705, -16, -256, -256, 15, -256, -256, -107, 164, -256, -256, 108, -256, -256),
                (-69, 126, -35, 491, -256, -256, -198, -256, -256, 698, -165, -256, -256, -146, -256, -256, 1133, 849, 220, -256, -256, 553, -256, -256, 757, 39, -256, -256, 1971, -256, -256),
                (885, 1053, 665, 220, -256, -256, 111, -256, -256, -143, 1054, -256, -256, 168, -256, -256, 473, 270, 325, -256, -256, 228, -256, -256, 2191, 1971, -256, -256, 298, -256, -256),
                (-71, 482, 496, 221, -256, -256, 472, -256, -256, 614, 91, -256, -256, 639, -256, -256, 109, 37, -26, -256, -256, 147, -256, -256, -107, 215, -256, -256, 381, -256, -256),
                (70, 83, 219, 147, -256, -256, -183, -256, -256, 733, 238, -256, -256, 35, -256, -256, 75, 271, 388, -256, -256, 2, -256, -256, 164, 1, -256, -256, -107, -256, -256),
                (218, -17, 327, 219, -256, -256, 383, -256, -256, 91, 73, -256, -256, 95, -256, -256, 207, 207, 513, -256, -256, 208, -256, -256, -67, -118, -256, -256, -36, -256, -256),
                (-30, 506, 350, 296, -256, -256, -262, -256, -256, -202, 4, -256, -256, -98, -256, -256, -159, -6, 338, -256, -256, -215, -256, -256, -21, 147, -256, -256, 62, -256, -256),
                (221, 205, 147, -71, -256, -256, -51, -256, -256, 420, 106, -256, -256, 427, -256, -256, 125, -183, -6, -256, -256, -6, -256, -256, 150, 822, -256, -256, -107, -256, -256),
                (494, 705, 452, 221, -256, -256, 104, -256, -256, -117, 1405, -256, -256, 226, -256, -256, 350, 676, -17, -256, -256, 216, -256, -256, 25, 634, -256, -256, 182, -256, -256),
                (1284, 1340, 1032, 220, -256, -256, 893, -256, -256, 289, 265, -256, -256, 140, -256, -256, 1337, 755, 754, -256, -256, 4328, -256, -256, 81, 1916, -256, -256, 1473, -256, -256),
                (-3, 200, -95, -35, -256, -256, 138, -256, -256, -201, -16, -256, -256, -16, -256, -256, -110, -6, 356, -256, -256, -159, -256, -256, 68, 586, -256, -256, 75, -256, -256),
                (494, 351, 615, -71, -256, -256, -53, -256, -256, 151, 243, -256, -256, 312, -256, -256, 174, 1618, 158, -256, -256, 747, -256, -256, -107, 263, -256, -256, 164, -256, -256),
                (885, 1053, 777, 221, -256, -256, 178, -256, -256, -185, 1054, -256, -256, 162, -256, -256, 482, 270, -53, -256, -256, 200, -256, -256, 2191, 2655, -256, -256, 915, -256, -256),
                (496, 705, 452, 220, -256, -256, 94, -256, -256, -142, 320, -256, -256, 226, -256, -256, 350, 676, -17, -256, -256, 216, -256, -256, 25, 634, -256, -256, 182, -256, -256),
                (349, 14, 147, -30, -256, -256, -17, -256, -256, 63, 115, -256, -256, 164, -256, -256, -13, 462, 73, -256, -256, -60, -256, -256, 639, 349, -256, -256, 86, -256, -256),
                (218, -36, -66, -202, -256, -256, 1, -256, -256, 377, -96, -256, -256, -17, -256, -256, 201, 513, 523, -256, -256, 543, -256, -256, 381, -77, -256, -256, 1141, -256, -256),
                (514, 351, 381, 302, -256, -256, 93, -256, -256, 151, 243, -256, -256, 312, -256, -256, 464, 676, 164, -256, -256, 216, -256, -256, 1108, 869, -256, -256, 787, -256, -256),
                (1536, 1032, 1412, 220, -256, -256, 1399, -256, -256, -35, 325, -256, -256, -16, -256, -256, 1785, 167, 1931, -256, -256, 266, -256, -256, 1795, 2410, -256, -256, 43, -256, -256),
                (218, -35, 172, 200, -256, -256, 222, -256, -256, 91, 73, -256, -256, -84, -256, -256, 201, 197, 1204, -256, -256, 103, -256, -256, 381, -77, -256, -256, -49, -256, -256),
                (-63, 126, -35, 491, -256, -256, -197, -256, -256, 748, -165, -256, -256, -236, -256, -256, 849, 665, 220, -256, -256, 89, -256, -256, 607, 322, -256, -256, 279, -256, -256),
                (220, 215, 147, -89, -256, -256, -18, -256, -256, 200, -17, -256, -256, 340, -256, -256, 108, -159, -6, -256, -256, 430, -256, -256, 164, 115, -256, -256, -67, -256, -256),
                (19, 186, -60, -35, -256, -256, 98, -256, -256, -201, -16, -256, -256, -16, -256, -256, 68, 259, -193, -256, -256, 586, -256, -256, 62, 91, -256, -256, 164, -256, -256),
                (494, 351, 452, -71, -256, -256, 405, -256, -256, -259, 383, -256, -256, -6, -256, -256, 174, 2078, 158, -256, -256, 747, -256, -256, -53, 2750, -256, -256, 164, -256, -256),
                (200, -114, 4, 351, -256, -256, -215, -256, -256, 851, 899, -256, -256, 622, -256, -256, 462, 210, -67, -256, -256, -67, -256, -256, 886, -45, -256, -256, 190, -256, -256),
                (334, 348, 615, -30, -256, -256, 172, -256, -256, 99, -259, -256, -256, 658, -256, -256, 166, 127, 383, -256, -256, 357, -256, -256, -53, 263, -256, -256, 164, -256, -256),
                (514, 537, 482, 222, -256, -256, 115, -256, -256, -61, -211, -256, -256, 228, -256, -256, 196, 208, 197, -256, -256, 1826, -256, -256, -125, 158, -256, -256, 513, -256, -256),
                (1272, 1052, 44, 147, -256, -256, 62, -256, -256, 244, 538, -256, -256, 768, -256, -256, 1785, 289, 76, -256, -256, 2582, -256, -256, 31, -9, -256, -256, 4404, -256, -256),
                (484, 659, 452, 221, -256, -256, 94, -256, -256, 65, 1, -256, -256, 126, -256, -256, 145, 567, 109, -256, -256, 816, -256, -256, 676, -67, -256, -256, 828, -256, -256),
                (265, 70, 56, 199, -256, -256, -176, -256, -256, 63, 752, -256, -256, 164, -256, -256, 91, 55, 377, -256, -256, 1138, -256, -256, 482, 164, -256, -256, 145, -256, -256),
                (334, 356, 615, -40, -256, -256, -53, -256, -256, 158, -259, -256, -256, 1123, -256, -256, 391, 93, 15, -256, -256, -17, -256, -256, 440, 80, -256, -256, 193, -256, -256),
                (218, -121, -16, 103, -256, -256, -199, -256, -256, 851, 899, -256, -256, 622, -256, -256, 201, 513, 523, -256, -256, 543, -256, -256, 238, -36, -256, -256, -49, -256, -256),
                (-3, 105, -95, -35, -256, -256, -66, -256, -256, -172, -77, -256, -256, 317, -256, -256, 5, 147, 221, -256, -256, 157, -256, -256, 62, 91, -256, -256, 164, -256, -256),
                (334, 356, 615, -53, -256, -256, -53, -256, -256, 158, 130, -256, -256, 1123, -256, -256, 166, 1618, 127, -256, -256, -169, -256, -256, -53, 263, -256, -256, 164, -256, -256),
                (885, 821, 1184, 1164, -256, -256, 289, -256, -256, 25, -26, -256, -256, 155, -256, -256, 270, 325, 238, -256, -256, 340, -256, -256, -17, 887, -256, -256, 3, -256, -256),
                (250, 356, 360, 220, -256, -256, 93, -256, -256, 83, -242, -256, -256, 387, -256, -256, 115, 25, 48, -256, -256, 391, -256, -256, -35, 125, -256, -256, 164, -256, -256),
                (109, 1, 167, 197, -256, -256, -26, -256, -256, 181, -23, -256, -256, 68, -256, -256, -97, 242, 182, -256, -256, 249, -256, -256, -67, 222, -256, -256, -246, -256, -256),
                (334, 554, 1113, 482, -256, -256, 182, -256, -256, -80, 1405, -256, -256, 91, -256, -256, 166, 165, 391, -256, -256, 767, -256, -256, -53, 86, -256, -256, 164, -256, -256),
                (265, 70, 147, -30, -256, -256, -17, -256, -256, 63, 752, -256, -256, 164, -256, -256, 91, 55, 117, -256, -256, 1138, -256, -256, 482, 164, -256, -256, 145, -256, -256),
                (482, 659, 452, 221, -256, -256, -39, -256, -256, -50, -36, -256, -256, 1479, -256, -256, 309, 218, 220, -256, -256, 162, -256, -256, 25, 634, -256, -256, 55, -256, -256),
                (1272, 849, 103, 147, -256, -256, 115, -256, -256, 745, 229, -256, -256, 146, -256, -256, 1785, 289, 359, -256, -256, 73, -256, -256, 31, -9, -256, -256, 1298, -256, -256),
                (263, 356, -23, 147, -256, -256, 220, -256, -256, 115, -107, -256, -256, 402, -256, -256, 167, 127, 55, -256, -256, -107, -256, -256, -35, 167, -256, -256, 258, -256, -256),
                (152, 221, -35, 289, -256, -256, 109, -256, -256, -122, -6, -256, -256, 46, -256, -256, 115, 822, 238, -256, -256, 258, -256, -256, -35, 123, -256, -256, 164, -256, -256)
                );
    constant value_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 0, 0, 0, 386, -11, 0, 1, 21, 2, 1, 115, 35, 3, 80, 126, 6, 5, 7, 174, 302, 4, 106, 175, 9, 8, 285, 228, 10, 320, 241),
                (0, 0, 0, 0, 31, -11, 0, -4, 9, 1, 1, 38, 13, 2, 27, 43, 4, 3, 2, 59, 34, 4, 45, 34, 6, 7, 40, 45, 5, 44, 37),
                (0, 0, 0, 0, 27, -11, 0, -4, 8, 1, 0, 23, 7, 1, 19, 29, 4, 3, 2, 33, 23, 4, 33, 25, 5, 6, 29, 34, 4, 30, 28),
                (0, 0, 0, 24, 0, -11, -4, 1, 0, 4, 14, 1, 27, 14, 3, 2, 3, 31, 12, 2, 13, 20, 4, 5, 24, 28, 4, 22, 23, 24, 24),
                (0, 0, 0, 0, 22, -11, 0, -5, 4, 1, 0, 6, 16, 1, 20, 4, 3, 2, 5, 27, 31, 2, 12, 17, 4, 5, 20, 24, 3, 18, 19),
                (0, 0, 0, 21, 0, -11, -5, 0, 0, 8, -1, 1, 14, 3, 3, 2, 2, 20, 10, 1, 7, 13, 4, 4, 17, 21, 3, 14, 17, 21, 21),
                (0, 0, 0, 20, 0, -10, -1, 0, 0, 8, -1, 1, 15, 4, 2, 1, 4, 18, 25, 1, 8, 12, 3, 4, 15, 19, 3, 12, 14, 20, 20),
                (0, 0, 0, 19, 0, -10, -2, 0, 0, 14, 3, 1, 12, 2, 2, 1, 4, 15, 22, 1, 7, 10, 3, 3, 13, 18, 2, 10, 13, 19, 19),
                (0, 0, 0, 18, 0, -11, -5, 0, 0, 8, 0, 1, 5, 9, 2, 1, 1, 10, 1, 2, 19, 8, 3, 3, 13, 17, 2, 12, 3, 18, 18),
                (0, 0, 0, 17, 0, -1, -9, 0, 0, 2, 18, 0, -3, 4, 2, 1, 3, 13, 17, 1, 5, 8, 3, 3, 12, 15, 2, 11, 4, 17, 17),
                (0, 0, 0, 0, 17, -10, 0, 17, -2, 0, 0, 15, 4, 0, -4, 3, 2, 1, 1, 11, 4, 1, 3, 5, 2, 3, 10, 14, 2, 7, 9),
                (0, 0, 0, 0, 16, 0, 0, -10, -3, 0, 0, 5, -3, 0, 17, 4, 1, 1, 1, 5, 12, 0, -1, 5, 2, 2, 9, 13, 2, 8, 1),
                (0, 0, 0, 3, 16, 16, 0, -1, -9, 0, 0, 0, 13, 0, 3, -3, 1, 1, 1, 11, 2, 1, 8, 3, 2, 2, 8, 12, 1, 4, 7),
                (0, 0, 0, 0, 16, -9, 0, 9, -1, 0, 0, 7, 14, 0, 18, -2, 1, 1, 1, 9, 3, 0, 2, 4, 2, 2, 11, 7, 1, 16, 6),
                (0, 0, 0, 0, 8, -7, 0, -8, -2, 0, 0, 13, 1, 1, 9, 0, 1, 1, 2, 7, 12, 1, 2, 5, 2, 2, 7, 10, 1, 6, 0),
                (0, 0, 0, 0, 2, 29, 0, -10, -4, 0, 0, 0, 11, 0, -5, -1, 1, 1, 1, 3, 9, 0, -3, 3, 1, 2, 7, 13, 1, -3, 6),
                (0, 0, 0, 2, 15, 16, 0, 0, -8, 0, 0, 8, 1, 1, 19, 10, 1, 1, 1, 6, 2, 0, 5, 1, 1, 1, 5, 8, 1, 5, -2),
                (0, 0, 0, 0, 6, -7, 0, 4, -4, 0, 1, 7, 1, 0, 2, 11, 1, 2, 3, 18, 16, 2, -4, 12, 1, 0, 3, -7, 1, 10, 4),
                (0, 0, 0, 0, 15, -8, 0, 9, 0, 0, 1, 6, 1, 0, 4, 1, 1, 1, 1, 3, 8, 1, -1, 4, 2, 2, 9, 13, -1, 5, -14),
                (0, 0, 0, 0, 1, -7, 0, 3, -5, 0, 0, 1, 6, 0, -4, 1, 1, 2, 3, 16, 15, 2, -4, 11, 1, 0, 4, -4, 1, 8, 3),
                (0, 0, 0, 0, 15, -8, 0, 8, -1, 0, 0, 1, 7, 0, 0, 8, 1, 1, 1, 2, 4, -1, 11, -9, 2, 2, -8, 9, -1, -7, 18),
                (0, 0, 0, 0, -7, -2, 0, 6, -3, 0, 0, 1, 7, 0, -4, 1, 1, 2, 2, 14, 12, 2, 8, 12, 1, 0, 2, -6, 1, 9, 3),
                (0, 0, 0, 0, 14, -6, 0, 8, -6, 0, 0, 1, 9, 0, -1, -2, 1, 1, 1, 4, 1, -1, 9, -10, 1, 1, 6, 9, 0, -7, 9),
                (0, 0, 0, 0, 10, -7, 0, -2, 3, 0, 0, 1, 4, 0, -1, -6, 1, 0, 2, 2, 8, 0, 3, -1, 1, 1, 7, 4, 0, -7, 5),
                (0, 0, 0, 0, 2, -7, 0, 11, 0, 0, 0, 1, 5, 0, -1, -12, 1, 1, 1, 5, 2, -2, 6, -12, 1, 1, 7, 11, 0, 12, -5),
                (0, 0, 0, 0, 12, -6, 0, 2, -3, 0, 0, 1, 5, 0, 0, -8, 0, 0, 1, 5, -3, 0, 1, -9, 1, 1, 3, 8, 0, -8, 7),
                (0, 0, 0, 0, 15, -6, 0, -2, 2, 0, 0, 0, 3, 0, -1, -10, 0, 0, 0, 4, 1, -1, 3, -6, 1, 1, 6, 14, -1, -13, 5),
                (0, 0, 0, 0, 7, -7, 1, 8, 2, 0, 0, -4, -4, 0, 7, 1, 0, 0, 1, 4, -3, 0, 1, -8, 1, 1, 2, 4, 0, -7, 6),
                (0, 0, 0, 0, 11, -8, 1, 12, 7, 0, 0, -3, -2, 0, 5, 0, 0, 1, 1, 5, 7, 0, 7, -4, 0, 0, 1, -8, 1, 4, 2),
                (0, 0, 0, 0, 3, 8, 3, 13, 17, 0, 0, -2, 2, 0, -6, -1, 0, 1, 1, 1, 6, 0, 7, -3, 0, 0, 1, -8, 0, 6, 2),
                (0, 0, 0, 0, -3, 8, 0, -7, -1, 0, 0, 1, 5, 0, 0, -8, 0, 0, 0, 3, -1, 0, 0, 6, 2, 1, 21, 5, 3, 3, 17),
                (0, 0, 0, 0, 1, 8, 1, 5, 10, 0, 0, -6, 1, -1, -5, -2, 0, 1, 0, 5, 0, 1, 5, 2, 0, 0, 0, -6, 0, 5, 2),
                (0, 0, 0, 0, -4, 5, 0, 2, -5, 0, 0, 5, 6, 0, -3, -3, 0, 1, 1, 1, 4, 0, 3, -5, 0, 0, 0, 4, 1, 21, 8),
                (0, 0, 0, 1, 14, 16, 0, 3, -5, 0, 0, 0, 5, 0, -1, -1, 0, 0, 0, 1, -5, 0, 6, 1, -1, -2, 5, -9, 1, 7, -4),
                (0, 0, 0, 0, 1, 7, 1, 4, 7, 0, 0, -1, 4, -2, -5, -12, 0, 0, 0, 2, 1, -1, -10, 0, 1, 2, 15, 22, 1, -3, 10),
                (0, 0, 0, 0, -6, 0, 0, 3, -1, 0, 1, -4, 5, 0, -5, -1, 0, 1, 0, 6, 1, 1, 6, 1, 0, 0, 0, 3, 0, 15, 5),
                (0, 0, 0, 0, 4, -4, 2, 12, 7, 0, 0, -5, 0, -1, -7, -2, 0, 1, 0, 7, 0, 1, 5, 1, 0, 0, 1, 5, 0, -3, 1),
                (0, 0, 0, 0, 2, -4, 0, 0, -5, 1, 1, 8, 10, -1, -15, -3, 0, 1, 0, 5, -3, 1, 10, 4, 0, 0, -1, 3, 0, 0, 5),
                (0, 0, 1, 1, 14, 14, 2, 15, 16, 0, 0, 4, -6, 0, 7, -1, 0, 0, 0, 5, 0, 1, 13, 4, 0, 0, -1, -2, 0, 5, 0),
                (0, 0, 0, 0, 6, -6, 1, 13, 7, 0, 0, 1, -5, 0, 1, -4, 0, 1, 0, 6, -2, 1, 9, 4, 0, 0, 1, 4, 0, 0, 1),
                (0, 0, 0, 0, 2, -4, 0, 1, -4, 1, 1, 7, 8, -2, -52, -6, 0, 1, 0, 5, -3, 1, 8, 4, 0, 0, 0, 4, 0, 0, 6),
                (0, 0, 0, 0, 1, -2, 1, 6, 1, -1, 1, 9, 2, -1, -9, -2, 0, 0, 0, 12, -2, 1, 4, 14, 0, 0, -41, 2, -2, -13, 2),
                (0, 0, 1, 1, 13, 14, 2, 15, 16, 0, 0, -8, 14, 0, -4, 10, 0, 0, 0, 0, 1, 0, 10, 2, 0, 0, 1, 7, 0, -4, 0),
                (0, 0, 0, 0, 5, -6, 1, 10, 5, 0, 0, 1, -5, -1, 0, -5, 0, 1, 0, 7, -1, 1, 8, 1, 0, 0, 3, 3, 0, 0, -3),
                (0, 0, 0, 0, 0, -1, 1, 5, 1, -1, 1, 5, -70, -1, -8, -2, 0, 0, 1, 15, 5, 0, -2, -30, 0, 1, 4, 7, 0, 3, -7),
                (0, 0, 0, 0, -2, 5, 0, 2, -3, 0, 0, 1, -5, 1, 3, 13, 0, 0, 0, -1, 10, 0, 6, 0, 0, 0, 3, 6, 0, -3, -1),
                (0, 0, 1, 1, 13, 14, 2, 14, 15, 0, 0, -6, 105, 0, 5, -4, 0, 0, 0, 3, -1, 0, 9, 2, 0, 0, 0, -3, 1, 6, -24),
                (0, 0, 0, 0, 0, -1, 0, 3, -2, -1, 0, 0, 7, -1, -11, -2, 0, 0, 0, 13, -9, 1, 66, 199, 1, 11, 314, 34, 1, 5, 11),
                (0, 0, 0, 0, -2, 1, 0, 3, 9, 0, 0, -2, 0, -1, -6, -2, 0, 0, 0, 3, -3, 0, 5, 1, -1, -1, 3, -8, 1, 5, -3),
                (0, 0, 0, 0, 1, -4, 0, 1, -4, 0, 1, 4, 9, -4, -53, -12, 0, 1, 0, 5, -2, 1, 7, -2, 0, 0, 2, 3, 0, 0, 4),
                (0, 0, 0, 0, -2, 4, 0, 2, -3, 0, 0, 1, -6, 1, 4, 15, 0, 0, 0, -1, 8, 0, 5, 0, 0, 0, 6, 10, 0, -1, 1),
                (0, 0, 0, 0, 14, -3, 0, 2, -1, 0, 0, 3, -1, 2, 21, 6, 0, 0, 0, -6, -2, -3, -28, -3, 0, 1, 4, 8, 0, -2, 0),
                (0, 0, 0, 0, 0, -1, 0, 2, -3, -1, 0, -2, 5, -2, -8, 23, 0, 0, 0, 11, -1, 1, 4, 11, -1, -3, 10, -17, 0, 3, -27),
                (0, 0, 0, 0, -1, -1, 0, 6, 1, 0, 1, 2, 8, -1, -10, -1, 0, 0, 0, 2, -4, 0, 24, 9, 0, 0, 2, 5, 0, -4, 0),
                (0, 0, 0, 0, 0, -1, 0, 4, 0, 0, 1, 15, 5, -1, -6, -1, 0, 0, -1, 9, -26, 0, 3, 16, -1, 1, -52, 7, -1, -18, -3),
                (0, 0, 0, 0, 1, -5, 0, -1, -7, 1, 1, 6, 12, -1, 5, -19, 0, 0, 0, 5, -3, 1, 6, 3, 0, 0, 1, 3, 0, -4, 0),
                (0, 0, 0, 0, -1, 2, 0, 4, -2, 0, 0, -2, 3, 0, -1, 2, 0, 0, 0, 275, 5, 0, 218, 20, 1, 1, 9, 14, 0, -5, 11),
                (0, 0, 0, 0, -1, -1, 0, 4, 1, 0, 0, 1, 9, 0, 7, -1, 0, 0, 0, -5, 52, 8, 71, -14, 0, -2, 4, -14, 0, 10, -3),
                (0, 0, 0, 0, 14, -3, 0, 1, 4, 0, 0, 3, -1, 1, 9, 3, 0, 0, 0, -3, -1, -3, -22, -2, 0, 1, 4, 7, 0, -1, 0),
                (0, 0, 0, 0, 0, 4, 0, 4, 2, 1, 1, 10, 5, 0, 4, -3, 0, 0, 0, 0, -1, 0, 1, 4, 0, -2, -6, -13, 0, 2, -3),
                (0, 0, 0, 0, 0, -1, 0, 3, 0, -1, 0, -51, 3, -1, -5, -16, 0, -1, -3, -1, -22, 0, -2, -14, 0, 0, 3, -1, -1, -5, 14),
                (0, 0, 0, 0, -2, -1, 0, 2, -19, 0, 1, 5, 2, 0, -4, 3, 0, 0, 0, 4, -1, 0, 2, 4, 0, 0, 2, 4, 0, -2, 1),
                (0, 0, 0, 0, 0, 5, 0, 1, -3, 0, 0, 1, 3, 0, 6, -2, 0, 0, 0, -1, 16, 0, 6, 8, 0, 0, 0, -3, 0, 27, 2),
                (0, 0, 0, 0, -1, -1, 0, 2, 0, 0, 0, 2, 7, 0, 0, -2, 0, 0, 0, -5, 13, 7, 47, -14, 0, -2, 3, -12, 0, 15, -2),
                (0, 0, 0, 0, -2, 2, -1, 1, -6, 0, 0, 3, 8, -4, 29, -19, 0, 0, 0, 4, -2, 1, 9, 4, 0, 0, 2, 2, 0, 1, 0),
                (0, 0, 0, 0, 1, -1, 0, 12, 1, 0, 0, 2, -1, 1, 17, 4, 0, 0, 0, -1, 6, 0, -5, -2, 0, 0, 1, -1, 0, 2, -2),
                (0, 0, 0, 0, 0, -1, 0, 3, -1, 0, 0, 3, -4, -1, -9, -3, 0, 0, 0, 2, -1, -1, 5, -9, 0, 1, 6, 4, 0, 0, 4),
                (0, 0, 0, 0, 0, 0, 0, 2, -2, -1, 0, -3, 5, -1, -5, -16, 0, 0, 0, 0, -144, 1, 4, 14, -1, -4, -24, -4, 0, 7, -3),
                (0, 0, 0, 0, 0, 7, 0, -4, -5, 0, 0, -1, 7, -1, -9, -3, 0, 0, 0, 3, -3, 1, 5, 2, 0, 0, 1, -2, 0, 1, -1),
                (0, 0, 0, 0, -1, 1, 0, 6, 0, 0, 0, -1, 1, -1, -8, -2, 0, 0, 0, 22, 2, -1, 0, -6, 0, 1, 5, 3, 0, -2, 3),
                (0, 0, 0, 0, 0, 0, 0, 2, -1, -1, 1, -33, 5, -1, -4, -14, 0, 0, -3, -3, -20, 0, -2, -20, 0, 0, 2, 7, -1, -20, -2),
                (0, 0, 0, 0, 0, -1, 0, 3, 0, 0, 0, 2, 8, -1, -7, -3, 0, 0, 0, 2, -1, -1, 4, -7, 0, 0, 6, 3, 0, 0, 3),
                (0, 0, 0, 0, -1, 1, 0, 0, 3, 0, 0, -2, 3, 0, -1, 2, 0, 0, 0, 9, -9, 2, 548, 40, 0, 1, 33, 6, 0, -5, 7),
                (0, 0, 0, 1, 13, 15, 0, -5, 0, 0, 0, 1, 0, 1, 12, 4, 0, 0, 0, -4, -17, 1, 62, 1, 0, -1, -9, -2, 0, 2, -6),
                (0, 0, 0, 0, 0, 5, 0, 4, 0, 0, 0, -1, 1, -1, -7, -1, 0, 0, 0, 0, 4, -1, 4, -4, 0, 0, 2, 4, 0, -4, 0),
                (0, 0, 0, 0, 0, 0, 0, 4, 11, 0, 1, 10, 3, 0, 17, 0, 0, -1, 0, -1, 13, -1, -16, -5, 0, 5, 17, 28, 0, -8, 3),
                (0, 0, 0, 0, -1, -1, 0, 0, 3, 0, 0, 1, 6, 0, 5, -1, 0, 0, 0, -4, 35, 1, 13, -11, 0, -1, -8, -2, 0, 9, 1),
                (0, 0, 0, 0, 0, 3, 0, 3, 2, 0, 1, 8, 3, 0, 14, -1, 0, 0, 0, 0, 0, 0, 3, 1, 0, -1, -10, -5, 0, 4, -1),
                (0, 0, 0, 0, -2, 0, 0, 7, 1, 0, 1, 1, 5, 0, -5, 15, 0, 0, 0, -1, 4, 0, -2, -5, 0, 0, 1, -1, 0, -9, 2),
                (0, 0, 0, 0, 0, 5, 0, -3, -3, 0, 0, 0, 6, -1, -7, -3, 0, 0, 0, 4, 1, 0, 3, -1, 0, 0, 3, -5, 0, -1, 2),
                (0, 0, 0, 0, -1, 1, 0, 2, -5, 0, 0, -2, 4, 0, -5, 0, 0, 0, 0, 19, 2, -1, 1, -8, 0, 0, 2, 13, 0, -2, 2),
                (0, 0, 0, 0, 1, -2, 0, 7, 3, 0, 0, 0, 2, 0, -5, 1, 0, 0, 0, -7, 0, 0, -6, -1, 0, 1, 20, 3, -1, -5, 13),
                (0, 0, 0, 0, -1, 1, 0, 4, 0, 0, 0, 3, -1, -1, -3, -12, 0, 0, 0, 2, 0, 0, 5, 2, 0, 0, 3, 1, 0, -2, 1),
                (0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 4, 0, -1, -6, -1, 0, 0, 3, 6, 24, 0, 1, -3, 0, 1, 10, 3, 0, -2, 1),
                (0, 0, 0, 0, 0, 1, 0, 0, -1, 0, 0, 5, 1, 0, -4, 4, 0, -1, 0, 6, -1, -1, -4, -10, 0, -1, 13, -22, 0, 3, 10),
                (0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 4, -10, -1, -2, -9, 0, 0, 0, 0, -6, 0, 3, 0, 0, 1, -6, 4, 0, -2, 2),
                (0, 0, 0, 0, 0, -1, 0, 5, 1, 0, 0, -1, 57, 0, -1, 2, 0, 0, 0, 2, 8, 0, 9, -18, 0, 0, -8, 4, -1, -20, -5),
                (0, 0, 0, 0, -3, 0, 0, 4, 0, 0, 0, 3, -1, -1, -7, 3, 0, 0, 1, 0, 5, 0, 2, -1, 0, 0, -4, 0, 0, 1, -1),
                (0, 0, 0, 0, 2, -1, 0, 5, 3, 0, 0, 0, 2, 0, -4, 1, 0, 0, 0, -4, -17, 1, 38, 1, 0, -1, 1, -4, 0, 4, 0),
                (0, 0, 0, 0, 0, 8, 0, 15, -3, 0, 0, -1, 2, 0, -3, -9, 0, 0, 0, 2, -1, 0, 9, 1, 0, 0, 3, -4, 0, -1, 1),
                (0, 0, 0, 0, -1, 1, 0, 4, 0, 0, 0, -2, 0, -1, -6, 3, 0, 0, 0, 1, 2, -1, 14, -4, 0, 0, 3, 1, 0, -2, 1),
                (0, 0, 0, 0, 0, -7, 1, 3, -6, 0, 0, 6, 0, -1, -2, -6, 0, -2, 0, 21, -13, -3, -40, -8, 0, 1, -40, 8, 0, -8, 1),
                (0, 0, 0, 0, 0, -1, 0, 3, 0, 0, 0, 2, -1, -1, -1, -5, 0, 0, 0, 1, 3, 0, 1, -1, 0, 0, -2, 1, 0, -2, 2),
                (0, 0, 0, 0, -1, -1, 0, 3, 0, 0, 0, 5, 3, 0, 3, -1, 0, 0, 0, 4, -5, 1, 14, 4, 0, 0, -6, -8, 0, 7, 0),
                (0, 0, 0, 0, 0, 1, 1, 3, 17, 0, 0, 1, -7, -1, -6, -1, 0, 0, 0, 2, 0, 2, 10, -5, 0, 0, 0, 2, 0, -1, 1),
                (0, 0, 0, 0, -1, 1, 0, 0, 2, 0, 0, -1, 34, 0, -1, 1, 0, 0, 0, 2, 2, 0, 8, -14, 0, 0, -7, 3, -1, -18, -5),
                (0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 6, -1, -1, -4, 3, 0, 0, 0, 1, -3, 1, 19, 4, 0, 0, 4, 2, 0, -4, 0),
                (0, 0, 0, 0, 0, 3, 0, 0, -1, 0, 0, 1, -2, 1, 10, 3, 0, 0, 0, -2, 4, -1, -2, -6, 0, -1, 12, -18, 0, -13, 4),
                (0, 0, 0, 0, 1, 3, 0, -1, -1, 0, 0, 5, -1, -1, -1, -7, 0, 0, 0, 1, -1, 0, 14, 2, 0, 0, -12, 1, 0, -2, 0),
                (0, 0, 0, 0, -1, 3, 0, 3, -1, 0, 0, -1, 2, 0, -4, -1, 0, 0, 0, 0, 2, 0, -5, 0, 0, 0, -3, 1, 0, -1, 1)
                );
    constant children_left : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 29, 5, -1, -1, 8, 9, -1, -1, 12, -1, -1, 15, 16, 17, -1, -1, 20, -1, -1, 23, 24, -1, -1, 27, -1, -1, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 29, 5, -1, -1, 8, 9, -1, -1, 12, -1, -1, 15, 16, 17, -1, -1, 20, -1, -1, 23, 24, -1, -1, 27, -1, -1, -1, -1),
                (1, 2, 3, 29, 5, -1, -1, 8, 9, -1, -1, 12, -1, -1, 15, 16, 17, -1, -1, 20, -1, -1, 23, 24, -1, -1, 27, -1, -1, -1, -1),
                (1, 2, 3, 29, 5, -1, -1, 8, 9, -1, -1, 12, -1, -1, 15, 16, 17, -1, -1, 20, -1, -1, 23, 24, -1, -1, 27, -1, -1, -1, -1),
                (1, 2, 3, 29, 5, -1, -1, 8, 9, -1, -1, 12, -1, -1, 15, 16, 17, -1, -1, 20, -1, -1, 23, 24, -1, -1, 27, -1, -1, -1, -1),
                (1, 2, 3, 29, 5, -1, -1, 8, 9, -1, -1, 12, -1, -1, 15, 16, 17, -1, -1, 20, -1, -1, 23, 24, -1, -1, 27, -1, -1, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1),
                (1, 2, 3, 4, -1, -1, 7, -1, -1, 10, 11, -1, -1, 14, -1, -1, 17, 18, 19, -1, -1, 22, -1, -1, 25, 26, -1, -1, 29, -1, -1)
                );
    constant children_right : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (14, 7, 4, 30, 6, -1, -1, 11, 10, -1, -1, 13, -1, -1, 22, 19, 18, -1, -1, 21, -1, -1, 26, 25, -1, -1, 28, -1, -1, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (14, 7, 4, 30, 6, -1, -1, 11, 10, -1, -1, 13, -1, -1, 22, 19, 18, -1, -1, 21, -1, -1, 26, 25, -1, -1, 28, -1, -1, -1, -1),
                (14, 7, 4, 30, 6, -1, -1, 11, 10, -1, -1, 13, -1, -1, 22, 19, 18, -1, -1, 21, -1, -1, 26, 25, -1, -1, 28, -1, -1, -1, -1),
                (14, 7, 4, 30, 6, -1, -1, 11, 10, -1, -1, 13, -1, -1, 22, 19, 18, -1, -1, 21, -1, -1, 26, 25, -1, -1, 28, -1, -1, -1, -1),
                (14, 7, 4, 30, 6, -1, -1, 11, 10, -1, -1, 13, -1, -1, 22, 19, 18, -1, -1, 21, -1, -1, 26, 25, -1, -1, 28, -1, -1, -1, -1),
                (14, 7, 4, 30, 6, -1, -1, 11, 10, -1, -1, 13, -1, -1, 22, 19, 18, -1, -1, 21, -1, -1, 26, 25, -1, -1, 28, -1, -1, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1),
                (16, 9, 6, 5, -1, -1, 8, -1, -1, 13, 12, -1, -1, 15, -1, -1, 24, 21, 20, -1, -1, 23, -1, -1, 28, 27, -1, -1, 30, -1, -1)
                );
    constant parent : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 2, 4, 4, 1, 7, 8, 8, 7, 11, 11, 0, 14, 15, 16, 16, 15, 19, 19, 14, 22, 23, 23, 22, 26, 26, 3, 3),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 2, 4, 4, 1, 7, 8, 8, 7, 11, 11, 0, 14, 15, 16, 16, 15, 19, 19, 14, 22, 23, 23, 22, 26, 26, 3, 3),
                (-1, 0, 1, 2, 2, 4, 4, 1, 7, 8, 8, 7, 11, 11, 0, 14, 15, 16, 16, 15, 19, 19, 14, 22, 23, 23, 22, 26, 26, 3, 3),
                (-1, 0, 1, 2, 2, 4, 4, 1, 7, 8, 8, 7, 11, 11, 0, 14, 15, 16, 16, 15, 19, 19, 14, 22, 23, 23, 22, 26, 26, 3, 3),
                (-1, 0, 1, 2, 2, 4, 4, 1, 7, 8, 8, 7, 11, 11, 0, 14, 15, 16, 16, 15, 19, 19, 14, 22, 23, 23, 22, 26, 26, 3, 3),
                (-1, 0, 1, 2, 2, 4, 4, 1, 7, 8, 8, 7, 11, 11, 0, 14, 15, 16, 16, 15, 19, 19, 14, 22, 23, 23, 22, 26, 26, 3, 3),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28),
                (-1, 0, 1, 2, 3, 3, 2, 6, 6, 1, 9, 10, 10, 9, 13, 13, 0, 16, 17, 18, 18, 17, 21, 21, 16, 24, 25, 25, 24, 28, 28)
                );
    constant depth : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 4, 4),
                (0, 1, 2, 3, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 4, 4),
                (0, 1, 2, 3, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 4, 4),
                (0, 1, 2, 3, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 4, 4),
                (0, 1, 2, 3, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4),
                (0, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4, 1, 2, 3, 4, 4, 3, 4, 4, 2, 3, 4, 4, 3, 4, 4)
                );
    constant iLeaf : intArray2D(nTrees-1 downto 0)(nLeaves-1 downto 0) := ((4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (5, 6, 9, 10, 12, 13, 17, 18, 20, 21, 24, 25, 27, 28, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (5, 6, 9, 10, 12, 13, 17, 18, 20, 21, 24, 25, 27, 28, 29, 30),
                (5, 6, 9, 10, 12, 13, 17, 18, 20, 21, 24, 25, 27, 28, 29, 30),
                (5, 6, 9, 10, 12, 13, 17, 18, 20, 21, 24, 25, 27, 28, 29, 30),
                (5, 6, 9, 10, 12, 13, 17, 18, 20, 21, 24, 25, 27, 28, 29, 30),
                (5, 6, 9, 10, 12, 13, 17, 18, 20, 21, 24, 25, 27, 28, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30),
                (4, 5, 7, 8, 11, 12, 14, 15, 19, 20, 22, 23, 26, 27, 29, 30)
                );
    constant value : tyArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_tyArray2D(value_int);
      constant threshold : txArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_txArray2D(threshold_int);
end Arrays0;